LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;

ENTITY slave_SPI IS
PORT(
	CK, MOSI, nSS, SCK, RST_S : IN STD_LOGIC;
	MISO: OUT STD_LOGIC
	);
END slave_SPI;

ARCHITECTURE behavior OF slave_SPI IS

COMPONENT SPI IS
PORT(
	CK, MOSI, nSS, SCK, RST_S : IN STD_LOGIC;
	DOUT : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	A : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	DIN : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	MISO, RD, WR : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT memory is
PORT(
  	 clk, RD, WRn : in STD_LOGIC;
	 address : in STD_LOGIC_VECTOR(7 DOWNTO 0);
 	 data_in : in STD_LOGIC_VECTOR(15 DOWNTO 0);
 	 data_out : out STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END COMPONENT;

SIGNAL DOUT, DIN : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL RD, WR, WRn :  STD_LOGIC;
SIGNAL A : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN

WRn <= not WR;

mem : memory PORT MAP(CK, RD, WRn, A, DIN, DOUT);
spi1 :SPI PORT MAP(CK, MOSI, nSS, SCK, RST_S, DOUT, A, DIN, MISO, RD, WR);

END behavior;
