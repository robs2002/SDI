LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY microrom IS
PORT(
  address : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
  data_out : OUT STD_LOGIC_VECTOR(27 DOWNTO 0)
);
END microrom;

ARCHITECTURE Behavioral OF microrom IS

TYPE memory IS ARRAY(0 TO 15) OF STD_LOGIC_VECTOR(27 DOWNTO 0);

constant myrom : memory := (
0 =>  "0100000000000000000000000000" ,
1 =>  "0000000000000101010000000000" , 
2 =>  "0000100000000010101000000000" , 
3 =>  "0000101000000000000000000000" , 
4 =>  "0000111000000000000100000000" , 
5 =>  "0000110010000000000100000000" , 
6 =>  "0000000100000000000110000000" , 
7 =>  "0101000000100000000110001100" ,
8 =>  "0001010000000101010001100000" ,
9 =>  "0000100001000010101011010000" , 
10 => "0000101001010000000000100000" , 
11 => "1010111000001000000100100101" , 
12 => "0001010000000000000001100000" ,
13 => "0000000001000000000011010000" , 
14 => "0000000001010000000000100000" , 
15 => "1010000000001000000000100000" ) ;

BEGIN

data_out <= myrom(TO_INTEGER(UNSIGNED(address)));


END Behavioral;
