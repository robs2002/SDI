library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY fft_tb IS
   
end fft_tb;

ARCHITECTURE test OF fft_tb IS

COMPONENT fft IS
PORT(
	X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, W0, W1, W2, W3, W4, W5, W6, W7 : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
	Start, Clock, Reset : IN STD_LOGIC;
	Done : OUT STD_LOGIC;
	X0p, X1p, X2p, X3p, X4p, X5p, X6p, X7p, X8p, X9p, X10p, X11p, X12p, X13p, X14p, X15p: OUT STD_LOGIC_VECTOR (23 DOWNTO 0)
);
END COMPONENT;

SIGNAL X0_tb, X1_tb, X2_tb, X3_tb, X4_tb, X5_tb, X6_tb, X7_tb, X8_tb, X9_tb, X10_tb, X11_tb, X12_tb, X13_tb, X14_tb, X15_tb,
X0p_tb, X1p_tb, X2p_tb, X3p_tb, X4p_tb, X5p_tb, X6p_tb, X7p_tb, X8p_tb, X9p_tb, X10p_tb, X11p_tb, X12p_tb, X13p_tb, X14p_tb, X15p_tb,
W0_tb, W1_tb, W2_tb, W3_tb, W4_tb, W5_tb, W6_tb, W7_tb : STD_LOGIC_VECTOR (23 DOWNTO 0); 
SIGNAL Start_tb, Clock_tb, Reset_tb, Done_tb : STD_LOGIC;

BEGIN

PROCESS
BEGIN
Clock_tb <= '0';
wait for 5 ns;
Clock_tb <= '1';
wait for 5 ns;
END PROCESS;

Reset_tb <= '1', '0' after 10 ns; 
Start_tb <= '0', '1' after 40 ns, '0' after 50 ns; 
X0_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "011111111111111111111111" after 55 ns, "000000000000000000000000" after 65 ns;
X1_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X2_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X3_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X4_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X5_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X6_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X7_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X8_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X9_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X10_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X11_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X12_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X13_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X14_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
X15_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 55 ns, "000000000000000000000000" after 65 ns;
W0_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "011111111111111111111111" after 55 ns, "000000000000000000000000" after 65 ns,
                                      "011111111111111111111111" after 155 ns, "000000000000000000000000" after 165 ns,
                                      "011111111111111111111111" after 265 ns, "000000000000000000000000" after 275 ns,
                                      "011111111111111111111111" after 375 ns, "000000000000000000000000" after 385 ns;
W1_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "011101100100000000000000" after 375 ns, "110011110001000000000000" after 385 ns;
W2_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "010110101000000000000000" after 265 ns, "101001011000000000000000" after 275 ns,
                                      "010110101000000000000000" after 375 ns, "101001011000000000000000" after 385 ns;
W3_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "001100001111000000000000" after 375 ns, "100010011100000000000000" after 385 ns;
W4_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "000000000000000000000000" after 155 ns, "100000000000000000000000" after 165 ns,
                                      "000000000000000000000000" after 265 ns, "100000000000000000000000" after 275 ns,
                                      "000000000000000000000000" after 375 ns, "100000000000000000000000" after 385 ns;
W5_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "110011110001000000000000" after 375 ns, "100010011100000000000000" after 385 ns;
W6_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "101001011000000000000000" after 265 ns, "101001011000000000000000" after 275 ns,
                                      "101001011000000000000000" after 375 ns, "101001011000000000000000" after 385 ns;
W7_tb <= "UUUUUUUUUUUUUUUUUUUUUUUU" , "100010011100000000000000" after 375 ns, "110011110001000000000000" after 385 ns;

fft_tb: fft PORT MAP (X0_tb, X1_tb, X2_tb, X3_tb, X4_tb, X5_tb, X6_tb, X7_tb, X8_tb, X9_tb, X10_tb, X11_tb, X12_tb, X13_tb, X14_tb, X15_tb,
		      W0_tb, W1_tb, W2_tb, W3_tb, W4_tb, W5_tb, W6_tb, W7_tb, Start_tb, Clock_tb, Reset_tb, Done_tb, X0p_tb, X1p_tb, X2p_tb, 
		      X3p_tb, X4p_tb, X5p_tb, X6p_tb, X7p_tb, X8p_tb, X9p_tb, X10p_tb, X11p_tb, X12p_tb, X13p_tb, X14p_tb, X15p_tb);

END test;
