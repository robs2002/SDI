library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY round_tb IS

END round_tb;

ARCHITECTURE test OF round_tb IS

COMPONENT round IS
PORT( DATA_IN : IN STD_LOGIC_VECTOR(48 DOWNTO 0);
	Clock, Reset : IN STD_LOGIC;
      DATA_OUT : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
);
END COMPONENT;

SIGNAL clk_tb, rst_tb: STD_LOGIC;
SIGNAL a_s: STD_LOGIC_VECTOR(48 DOWNTO 0);
SIGNAL p_s: STD_LOGIC_VECTOR(23 DOWNTO 0);

BEGIN

PROCESS
BEGIN
clk_tb <= '0';
wait for 5 ns;
clk_tb <= '1';
wait for 5 ns;
END PROCESS;

process
begin
a_s <= "0010000000000000000000000100000000000000000000000";
wait for 50 ns;
a_s <= "1110101010101010101010101010101010101010101010101";
wait for 50 ns;
a_s <= "1111111111111111111111111111111111111111111111111";
wait for 50 ns;
a_s <= "0000000000000000000000000000000000000000000000000";
wait for 50 ns;
a_s <= "1110000000000100000000001110000000000100000000000";
wait for 50 ns;
a_s <= "1110000000000100000000001100000000000000000000000";
wait for 50 ns;
a_s <= "1110000000000100000000000100000000000000000000000";
wait;
end process;

rst_tb <= '1', '0' after 10 ns;

dut: round GENERIC MAP(24) PORT MAP (a_s, clk_tb, rst_tb, p_s);

END test;